`timescale 1ns / 1ps

//======================================================================
// Module: seg_display (���������)
// Description: 8λ8������ܶ�̬ɨ������ģ�顣
//              ����һ��32λ����ֵ��ÿ4λ����һ��Ҫ�ڶ�Ӧ�������
//              ��ʾ��ʮ�������� (0-F)��
//              �����ѡ(seg)��λѡ(an)�źš�
//              �ϸ���ѭ {g,f,e,d,c,b,a} �Ķ�ѡ����˳��
//======================================================================
module seg_display(
    // --- ģ��ӿ� ---
    input         clk,         // ����: 100MHz ϵͳʱ��
    input         rst_n,       // ����: ȫ�ָ�λ
    input  [31:0] data,        // ����: Ҫ��ʾ��8������ (data[3:0] ��Ӧ���ұߵĵ�0λ)
    
    output reg [6:0] seg,        // ���: 7���� (��ѡ)
    output reg [7:0] an          // ���: 8λ��������ѡ�� (λѡ)
);

    //---------------------------------------------------------
    // 1. �ڲ��źŶ���
    //---------------------------------------------------------
    
    // ɨ��ʱ�ӷ�Ƶ��/��������
    // ʹ��18λ��������ɨ��Ƶ�� = 100MHz / (2^18) �� 381Hz��
    // ���Ƶ���㹻�죬������ȫ�о�������˸��
    reg [17:0] clk_div;
    
    // ��ǰ����ɨ��������λ�� (0-7)��
    // ����ֱ���÷�Ƶ�������ĸ�3λ��Ϊɨ��ָ�롣
    wire [2:0] scan_pos = clk_div[17:15];
    
    // ��32λ���������У�ѡ���ĵ�ǰҪ��ʾ��4λ���֡�
    reg [3:0] digit_to_display;

    //---------------------------------------------------------
    // 2. ɨ��ʱ������
    //---------------------------------------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            clk_div <= 0;
        else
            clk_div <= clk_div + 1; // �������еļ�����
    end
    
    //---------------------------------------------------------
    // 3. ���������߼� (������߼�)
    //---------------------------------------------------------
    always @(*) begin
        // --- ����A: ����ѡ�� (MUX) ---
        // ���ݵ�ǰɨ���λ��(scan_pos)����32λ��data�����У�ѡ����Ӧ��4λ��
        case (scan_pos)
            3'd0: digit_to_display = data[3:0];   // ɨ�����ұ�(��0λ)�������
            3'd1: digit_to_display = data[7:4];   // ɨ���1λ�������
            3'd2: digit_to_display = data[11:8];  // ...
            3'd3: digit_to_display = data[15:12];
            3'd4: digit_to_display = data[19:16];
            3'd5: digit_to_display = data[23:20];
            3'd6: digit_to_display = data[27:24];
            3'd7: digit_to_display = data[31:28]; // ɨ�������(��7λ)�������
            default: digit_to_display = 4'hF;     // �����ϲ��ᷢ����Ĭ����ʾF (Ϩ��)
        endcase

        // --- ����B: λѡ���� ---
        // ���ݵ�ǰɨ���λ��(scan_pos)������λѡ�ź� an (�͵�ƽ��Ч)��
        // ��ȷ�������κ�һ��˲�䣬ֻ��һ��an���ǵ͵�ƽ����ֻ��һ������ܱ����
        case (scan_pos)
            3'd0: an = 8'b11111110; // �������ұ�(��0λ)�������
            3'd1: an = 8'b11111101; // �����1λ�������
            3'd2: an = 8'b11111011; // ...
            3'd3: an = 8'b11110111;
            3'd4: an = 8'b11101111;
            3'd5: an = 8'b11011111;
            3'd6: an = 8'b10111111;
            3'd7: an = 8'b01111111; // ���������(��7λ)�������
            default: an = 8'b11111111; // Ĭ��ȫ������
        endcase
        
        // --- ����C: ��ѡ���� (4λת7λ) ---
        // ��ѡ����4λ����(digit_to_display)������ɶ�Ӧ��7���롣
        // �������ϸ���ѭ 7'b{g, f, e, d, c, b, a} ��ʽ��0��1�硿����
        case (digit_to_display)
            4'd0: seg = 7'b1000000;
            4'd1: seg = 7'b1111001;
            4'd2: seg = 7'b0100100;
            4'd3: seg = 7'b0110000;
            4'd4: seg = 7'b0011001;
            4'd5: seg = 7'b0010010;
            4'd6: seg = 7'b0000010;
            4'd7: seg = 7'b1111000;
            4'd8: seg = 7'b0000000;
            4'd9: seg = 7'b0010000;
            4'ha: seg = 7'b0001000; // A
            4'hb: seg = 7'b0000011; // b
            4'hc: seg = 7'b1000110; // C
            4'hd: seg = 7'b0100001; // d
            4'he: seg = 7'b0000110; // E
            4'hf: seg = 7'b0001110; // F
            default: seg = 7'b1111111; // �������(������Ч����)��ȫ��
        endcase
    end
endmodule