`timescale 1ns / 1ps

//==============================================================
// Module: timer (����������)
//==============================================================
module timer(
    input         clk,             // ���룺ϵͳ��ʱ�� (100MHz)
    input         rst_n,           // ���룺��λ�ź�

    input         start_10s,       // ���룺"��ʼ10���ʱ"����
    output        done_10s,        // �����"10�뵽�ˣ�"����

    input         start_20s,       // ���룺"��ʼ20���ʱ"����
    output        done_20s         // �����"20�뵽�ˣ�"����
);

    //---------------------------------------------------------
    // 1. ���峣�� (Ŀ��ֵ)
    //---------------------------------------------------------
    parameter TARGET_10S = 30'd1_000_000_000;
    parameter TARGET_20S = 31'd2_000_000_000;
    
    //---------------------------------------------------------
    // 2. �ڲ����� (���ĺ��Ĳ���)
    //---------------------------------------------------------
    reg [29:0] counter_10s;        // 10�붨ʱ���ļ�����
    reg        is_running_10s;     // 10�붨ʱ���Ƿ������У�(��/��)
    
    reg [30:0] counter_20s;        // 20�붨ʱ���ļ�����
    reg        is_running_20s;     // 20�붨ʱ���Ƿ������У�(��/��)

    //---------------------------------------------------------
    // 3. �����߼� (�����ι���)
    //---------------------------------------------------------
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            // ��λʱ�������ж�������ʼ��
            counter_10s <= 0;
            is_running_10s <= 0; // 0 ����"��"
            counter_20s <= 0;
            is_running_20s <= 0;
        end
        else begin
            // --- 10�������߼� ---
            if (start_10s) begin              // ���"��ʼ"��ť������...
                is_running_10s <= 1;          // ...������״̬Ϊ"�ǣ���������"...
                counter_10s <= 0;             // ...���Ҽ�������0��ʼ��
            end 
            else if (counter_10s == TARGET_10S - 1) begin // ���������������...
                is_running_10s <= 0;          // ...������״̬Ϊ"����ֹͣ"...
                counter_10s <= 0;             // ...���Ҽ��������㡣
            end 
            else if (is_running_10s == 1) begin // ���״̬��"��������"...
                counter_10s <= counter_10s + 1; // ...��ô�������ͼ�һ��
            end

            // --- 20�������߼� (��������ȫһ��) ---
            if (start_20s) begin
                is_running_20s <= 1;
                counter_20s <= 0;
            end 
            else if (counter_20s == TARGET_20S - 1) begin
                is_running_20s <= 0;
                counter_20s <= 0;
            end 
            else if (is_running_20s == 1) begin
                counter_20s <= counter_20s + 1;
            end
        end
    end

    //---------------------------------------------------------
    // 4. ����ź�
    //---------------------------------------------------------
    // "���"�ź� = (��������ֵ == Ŀ��ֵ - 1)
    assign done_10s = (counter_10s == TARGET_10S - 1);
    assign done_20s = (counter_20s == TARGET_20S - 1);

endmodule